/*
 * @Author       : 中北大学-聂怀昊
 * @Date         : 2024-06-26 10:10:46
 * @LastEditTime : 2024-06-26 10:10:54
 * @FilePath     : \ysyx\ysyx-workbench\npc\vsrc\IDU\ysyx_23060191_DEC.v
 * @Description  : 指令译码模块
 * 
 * Copyright (c) 2024 by 873040830@qq.com, All Rights Reserved. 
 */
`include "/mnt/ysyx/ysyx-workbench/npc/vsrc/defines.v"

module ysyx_23060191_DEC (
    input  [`CPU_WIDTH-1:0] inst,

    output   
);

endmodule //ysyx_23060191_DECS